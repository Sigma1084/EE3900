RC circuit (before switching)

r1 1 2 1
r2 2 3 2 
v1 1 0 dc 1V
v2 3 0 dc 2V
c1 2 0 1u

*transient analysis 
.tran 100u 5u uic
*defining the run-time control functions
.control
run
*plotting output voltages
*if you want to show the plot, uncomment the below line
*plot v(2)
wrdata 2_output.dat v(2)
+ title "Voltage across capacitor"
.endc
